`default_nettype none
`timescale 1ns / 1ps

module top_level(

);

endmodule

`default_nettype wire